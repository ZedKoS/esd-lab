library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity ControlSystem is
  port (

  );
end entity;

architecture Behavior of ControlSystem is
begin
end architecture;
